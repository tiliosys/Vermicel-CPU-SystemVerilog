//
// SPDX-License-Identifier: CERN-OHL-W-2.0
// SPDX-FileCopyrightText: 2023 Guillaume Savaton <guillaume.savaton@tiliosys.fr>
//

`default_nettype none

package Verdata_pkg;

    typedef int unsigned  word_t;
    typedef int signed    signed_word_t;
    typedef bit[3:0]      wstrobe_t;
    typedef byte unsigned byte_t;

endpackage

