
package virgule_pkg;

    typedef int unsigned word_t;
    typedef int signed   signed_word_t;
    typedef bit[3:0]     wstrobe_t;

endpackage
