
// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.

package Types_pkg;

    typedef int unsigned word_t;
    typedef int signed   signed_word_t;
    typedef bit[3:0]     wstrobe_t;

endpackage

